
module system (
	clk_clk,
	reset_reset_n,
	custom_pio_0_conduit_end_parport);	

	input		clk_clk;
	input		reset_reset_n;
	inout	[7:0]	custom_pio_0_conduit_end_parport;
endmodule
