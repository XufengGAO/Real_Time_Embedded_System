
module system (
	clk_clk,
	custompio_0_conduit_end_parport,
	reset_reset_n);	

	input		clk_clk;
	inout	[7:0]	custompio_0_conduit_end_parport;
	input		reset_reset_n;
endmodule
